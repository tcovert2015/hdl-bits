`timescale 1ns/1ps

module top ( input in, output out);

   assign out - in;
   
endmodule // top
